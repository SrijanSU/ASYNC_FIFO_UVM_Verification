package fifo_pkg;
`include "uvm_pkg.sv"
`include "uvm_macros.svh"
`include "defines.sv"
`include "async_fifo_write_sequence_item.sv"
`include "async_fifo_read_sequence_item.sv"
`include "async_fifo_write_sequencer.sv"
`include "async_fifo_read_sequencer.sv"
`include "async_fifo_write_sequence.sv"
`include "async_fifo_read_sequence.sv"
`include "async_fifo_virtual_sequencer.sv"
`include "async_fifo_virtual_sequence.sv"
`include "async_fifo_write_driver.sv"
`include "async_fifo_read_driver.sv"
`include "async_fifo_write_monitor.sv"
`include "async_fifo_read_monitor.sv"
`include "async_fifo_write_agent.sv"
`include "async_fifo_read_agent.sv"
`include "async_fifo_scoreboard.sv"
`include "async_fifo_subscriber.sv"
`include "async_fifo_environment.sv"
`include "async_fifo_test.sv"
endpackage
