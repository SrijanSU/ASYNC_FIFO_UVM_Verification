`define DATA_WIDTH 8
`define ADDR_WIDTH 4
`define WRITE_CLK  5
`define READ_CLK   10

